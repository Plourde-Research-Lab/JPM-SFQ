* Inverter cell for AK library.  ak3tl201       Revised: Monday, April 25, 2016
* root                                          Revision: 6
* HYPRES, Inc.
*
*
*
*
P1 1 0 P1
Xdcsfq 1 2 dcsfq
XTL1 2 3 BJTL5
* XTL2 3 4 BJTL5
XOUT 3 stdout
.SUBCKT DCSFQ IN OUT
L1 IN N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
Lj1 N004530 N005070 L?
Lj2 N005071 0 L?
Lj3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 OUT JTL1
.ENDS
.SUBCKT JTL1  IN OUT
L1 IN N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 OUT L3*xl
J1 IN 0 J
J2 N002320 0 J(J1)
.SUBCKT BJTL IN OUT
L1 IN OUT L?
J1 OUT 0 JT(J1)
.ENDS
.SUBCKT BJTL5 IN OUT
XBJTL1 IN N1 BJTL
XBJTL2 N1 N2 BJTL
XBJTL3 N2 N3 BJTL
XBJTL4 N3 N4 BJTL
XBJTL5 N4 OUT BJTL
.ENDS
.SUBCKT stdout  IN
R1 N006161 0 0.5
L2 IN N006421 0.75*XL
L3 N006421 N005260 0.75*XL
I1 N006421 0 2.8*XI
L4 N005260 N005261 1.5*XL
I2 N005700 0 2.8*XI
L5 N005261 N005700 0.75*XL
L6 N005700 N005520 0.75*XL
L7 N005520 N006161 2*XL
J1 IN 0 J(2)
J2 N005260 0 J(2)
J3 N005261 0 J(2)
J4 N005520 0 J(2)
.ENDS
.END
