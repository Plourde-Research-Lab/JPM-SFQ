*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
P1 N00284 0 P1
XDCSFQ N00284 N50214 DCSFQ
XMSPL N50214 N00143 N00168 SPL1
XTL1 N00143 N00215 BJTL5
M1 0 llm(LC, LJ1, LM1)
LJ1   N00215 N01215 L1
J1   N01215 0      JT(J1)
XTL3 N01215 N00217 BJTL5
XBTL1 N00217 N00218 JTL1
XBTL2 N00218 N00219 JTL2
R1 N00219 0 R1
* P2 N10284 0 P1
* XDCSFQ2 N10284 N10214 DCSFQ
XTL21 N00168 N10215 BJTL5
M21 0 llm(LC, LJ21, -LM1)
LJ21   N10215 N61215 L1
J21   N61215 0     JT(J1)
XTL23 N61215 N10217 BJTL5
XBTL21 N10217 N10218 JTL1
XBTL22 N10218 N10219 JTL2
R2 N10219 0 R1
IC N20217 0 IC
LC N20217 0 LC
.SUBCKT DCSFQ IN OUT
L1 IN N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
Lj1 N004530 N005070 L?
Lj2 N005071 0 L?
Lj3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 OUT JTL0
.ENDS
.SUBCKT JTL0 IN OUT
L1 IN N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 OUT L3*xl
J1 IN 0 JJ
J2 N002320 0 JJ
.ENDS
.SUBCKT JTL1 IN OUT
L1 IN N002521 L1*xl
J1 N002521 0 J(J1)
L2 N002521 N003521 L1
L3 N003521 N002320 L1*xl
I1 N003521 0 I1*xi
L4 N002320 OUT L1*xl
J2 N002320 0 J(J1)
.ENDS
.SUBCKT JTL2 IN OUT
L1 IN N002521 L1*xl
J1 N002521 0 J(J1)
L2 N002521 N003521 L1
L3 N003521 N002320 L1*xl
I1 N003521 0 I1*xi
L4 N002320 OUT L1*xl
J2 N002320 0 J(J1)
.ENDS
.SUBCKT BJTL5 IN OUT
L1 IN N1 L1
J1 N1 0 JT(J1)
L2 N1 N2 L1
J2 N2 0 JT(J1)
L3 N2 N3 L1
I3 N3 0 I1
J3 N3 0 JT(J1)
L4 N3 N4 L1
J4 N4 0 JT(J1)
L5 N4 OUT L1
J5 OUT 0 JT(J1)
.ENDS
.SUBCKT SPL1 IN OUT1 OUT2
L1 N020660 N01976 L1*XL
L2 N01976 N021021 L1*XL
I1 N01976 0 I1*XI
L3 IN N01976 L1*XL
L4 OUT1 N020660 L2*XL
L5 N021021 OUT2 L2*XL
J1 N020660 0 JJ
J2 N021021 0 JJ
J3 IN 0 JJ
.ENDS
