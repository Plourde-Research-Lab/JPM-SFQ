*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
P1 1 0 P1
XMIN 1 2 stdin1
XT 2 3 TFF
XMOUT 3 stdout1
.SUBCKT TFF IN OUT
LJ2 N001321 N00332 LJ2
LJ3 N001641 0 LJ3
LJ5 N001801 0 LJ5
LJ4 N001481 N00316 LJ4
L1 N00332 N00475 L1
L2 N00475 OUT L2
I1 N000521 0 I1
L3 IN N000361 L3
L4 N000521 N00336 L4
L5 N000361 N000521 L5
J1 N000361 0 JJ
J2 N00336 N001321 JJ
J3 N00332 N001641 JJ
J4 N00336 N001481 JJ
J5 N00316 N001801 JJ
Lq1 N00475 N00316 Lq1
.ENDS
.SUBCKT STDOUT1  1
R1 N248211 0 0.5
L1 1 N24787 L1*xl
L2 N247991 N248211 2.0
XMT1 N24787 N247991 JTL
.ENDS
.SUBCKT JTL  1 2
L1 1 N003961 L1*xl
L2 N003961 2 L1*xl
I1 N003961 0 i1*xi
J1 1 0 J
J2 2 0 J(J1)
.ENDS
.SUBCKT STDIN1  1 2
L1 1 N00519 2
XM1 N00519 N00499 JTL1
XM2 N00499 2 JTL1
.ENDS
.SUBCKT JTL1  1 2
L1 1 N002781 L1*xl
L2 N002781 N002921 L1*xl
L3 N002921 2 L3*xl
I1 N002781 0 i1*xi
J1 1 0 J
J2 N002921 0 J(J1)
.ENDS
