* SFQ Qbit control                              Revised: Wednesday, February 21, 2018
* root                                          Revision: 2
* A.Kirichenko, HYPRES, INC.
* 
* 
* 
* 
L1 N093800 N093091 L1
L2 N093331 N094351 L2
I1 N056311 0 I1
I2 N09194 0 I2*XI2
I3 N09274 0 I3*XI3
C1 N093800 0 C1
C2 N094351 0 C2
XM1 N09052 N056311 dcsfq
XM3 N09246 N09134 N09052 SPL1
XM4 N09134 N090130 N09194 sw
XM5 N09246 N092120 N09274 sw
XMt1 N090130 N10199 jtl2
XPTL1   N10207 N093091 PTL10
XMt2 N092120 N10267 jtl2
XMt3 N10199 N10207 trx
XPTL2   N10259 N093331 PTL10
XMt4 N10267 N10259 trx
.SUBCKT trx  1 2
L1 1 N07575 ?
L2 N07575 N076091 L2*xl
I1 N07575 0 i?
J1 N07575 0 JJJ
Rq N076091 2 ?
.ENDS
.SUBCKT PTL10  1 2
XMACRO10   N002001 2 PTL
XMACRO1   1 N000481 PTL
XMACRO2   N000481 N000741 PTL
XMACRO3   N000741 N000921 PTL
XMACRO4   N000921 N001081 PTL
XMACRO5   N001081 N001281 PTL
XMACRO6   N001281 N001441 PTL
XMACRO7   N001441 N001641 PTL
XMACRO8   N001641 N001801 PTL
XMACRO9   N001801 N002001 PTL
.ENDS
.SUBCKT PTL  1 2
L1 1 N000561 L1
L2 N000561 N001301 L1
L3 N001301 N001891 L1
L4 N001891 N002361 L1
L5 N002361 N002841 L1
L6 N002841 N003331 L1
C1 N000561 0 C1
L7 N003331 N003831 L1
C2 N001301 0 C1
L8 N003831 N004331 L1
L9 N004331 N004840 L1
C3 N001891 0 C1
C4 N002361 0 C1
C5 N002841 0 C1
C6 N003331 0 C1
C7 N003831 0 C1
C8 N004331 0 C1
C9 N004840 0 C1
C10 2 0 C1
L10 N004840 2 L1
.ENDS
.SUBCKT jtl2  1 2
L0 1 N003400 L0*xl
L1 N003400 N003781 L1*xl
L2 N003781 N003200 L2*xl
L3 N003200 2 L3*xl
I1 N003781 0 i1*xi
J1 N003400 0 JJ
J2 N003200 0 JJ
.ENDS
.SUBCKT sw  1 2 3
Li1 3 N00861 0.1
L1 N007750 N00861 L1*xl
L2 N00861 N007891 L2*xl
L3 N007891 N00887 L3*xl
J1 N00825 N007750 JJ
J2 N007891 0 JJ
XM1 1 N00825 JTL
XM2 N00887 2 JTL
.ENDS
.SUBCKT JTL  1 2
L1 1 N006570 L1*xl
L2 N006570 2 L1*xl
I1 N006570 0 i1*xi
J1 1 0 J
J2 2 0 J(j1)
.ENDS
.SUBCKT SPL1  1 2 3
L1 N020660 N01976 L1*XL
L2 N01976 N021021 L1*XL
I1 N01976 0 I1*XI
L3 3 N01976 L1*XL
L4 1 N020660 L2*XL
L5 N021021 2 L2*XL
J1 N020660 0 JJ
J2 N021021 0 JJ
J3 3 0 JJ
.ENDS
.SUBCKT dcsfq  1 2
L1 2 N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
Lj1 N004530 N005070 L?
Lj2 N005071 0 L?
Lj3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 1 JTL1
.ENDS
.SUBCKT JTL1  1 2
L1 1 N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 2 L3*xl
J1 1 0 J
J2 N002320 0 J(J1)
.ENDS
.END
