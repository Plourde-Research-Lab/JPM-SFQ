* spice netlist for InductEx4 user manual example 5
* Inductors
LJPM      1   2   1000
*LJTLA     3   4   41
*LJTLB     5   6   41
LBias     7   8
KBias     LBias LJPM
* Ports
P1     1   2
*P2     3   4
*P3     5   6
P4     7   8
.end
