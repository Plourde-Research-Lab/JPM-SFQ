*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
IJPM N20217 0 IJPM*xi
LJPM N20217 0 LJPM*xl
P1 N00284 0 P1
XIN N00284 N50214 DCSFQ
XMSPL N50214 N00143 N00168 SPL1
XTL1 N00143 N00215 BJTL5
M1 0 llm(LJPM, LJ1, M1*xm)
LJ1   N00215 N01215 LJTL*xl
J1   N01215 0      JT(J1*xj)
XTL3 N01215 N00217 BJTL5
XBTL1 N00217 N00218 JTL1
* XBTL2 N00218 N00219 JTL2
XTL21 N00168 N10215 BJTL5
M21 0 llm(LJPM, LJ21, -M1*xm)
LJ21   N10215 N61215 LJTL*xl
J21   N61215 0     JT(J1*xj)
XTL23 N61215 N10217 BJTL5
XBTL21 N10217 N10218 JTL1
* XBTL22 N10218 N10219 JTL2
R1 N00218 0 R
R2 N10218 0 R
* XDFF N10219 N00219 N20219 DFF
* XOUT N20219 STDOUT
.SUBCKT DCSFQ IN OUT
L1 IN N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
Lj1 N004530 N005070 L?
Lj2 N005071 0 L?
Lj3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 OUT JTL0
.ENDS
.SUBCKT JTL0 IN OUT
L1 IN N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 OUT L3*xl
J1 IN 0 J(J1*xj)
J2 N002320 0 J(J1*xj)
.ENDS
.SUBCKT JTL1 IN OUT
L1 IN N002521 L1*xl
J1 N002521 0 J(J1*xj)
L2 N002521 N003521 L1
L3 N003521 N002320 L1*xl
I1 N003521 0 I1*xi
L4 N002320 OUT L1*xl
J2 N002320 0 J(J1*xj)
.ENDS
* .SUBCKT JTL2 IN OUT
* L1 IN N002521 L1*xl
* J1 N002521 0 J(J1)
* L2 N002521 N003521 L1
* L3 N003521 N002320 L1*xl
* I1 N003521 0 I1*xi
* L4 N002320 OUT L1*xl
* J2 N002320 0 J(J1)
* .ENDS
.SUBCKT JTL2 IN OUT
L1 IN N002521 L1*xl
J1 N002521 0 J(J1*xj)
L2 N002521 N003521 L1*xl
L3 N003521 OUT L1*xl
I1 N003521 0 I1*xi
J2 OUT 0 J(J1*xj)
.ENDS
.SUBCKT SPL1 IN OUT1 OUT2
L1 N020660 N01976 L1*XL
L2 N01976 N021021 L1*XL
I1 N01976 0 I1*XI
L3 IN N01976 L1*XL
L4 OUT1 N020660 L2*XL
L5 N021021 OUT2 L2*XL
J1 N020660 0 J(J1*xj)
J2 N021021 0 J(J2*xj)
J3 IN 0 J(J3*xj)
.ENDS
.SUBCKT TFF IN OUT
LJ2 N001321 N00332 LJ2
LJ3 N001641 0 LJ3
LJ5 N001801 0 LJ5
LJ4 N001481 N00316 LJ4
L1 N00332 N00475 L1
L2 N00475 OUT L2
I1 N000521 0 I1
L3 IN N000361 L3
L4 N000521 N00336 L4
L5 N000361 N000521 L5
J1 N000361 0 JJ
J2 N00336 N001321 JJ
J3 N00332 N001641 JJ
J4 N00336 N001481 JJ
J5 N00316 N001801 JJ
Lq1 N00475 N00316 Lq1
.ENDS
.SUBCKT JTL IN OUT
L1 IN N00487 L1*xl
L2 N00487 N00407 L1*xl
I1 N00407 0 I1*xi
L3 N00407 N00507 L1*xl
L4 N00507 OUT L1*xl
J1 N00487 0 J(J1*xj)
J2 N00507 0 J(J1*xj)
.ENDS
.SUBCKT DFF CLK IN OUT
LJ1 CLK N008111 LJ1
L1 IN N006930 L1
L2 N006930 OUT L2
Lj2 N007211 0 LJ2
J1 N008111 N006930 JJ
J2 OUT N007211 JJ
.ENDS
.SUBCKT BJTL5 IN OUT
L1 IN N1 L1*xl
J1 N1 0 JT(J1*xj)
L2 N1 N2 L1*xl
J2 N2 0 JT(J1*xj)
L3 N2 N3 L1*xl
J3 N3 0 JT(J1*xj)
L4 N3 OUT L1*xl
J4 OUT 0 JT(J1*xj)
* L5 N4 OUT L1*xl
* J5 OUT 0 JT(J1*xj)
.ENDS
.SUBCKT stdout IN
R1 N006161 0 0.5
L2 IN N006421 0.75*XL
L3 N006421 N005260 0.75*XL
I1 N006421 0 2.8*XI
L4 N005260 N005261 1.5*XL
I2 N005700 0 2.8*XI
L5 N005261 N005700 0.75*XL
L6 N005700 N005520 0.75*XL
L7 N005520 N006161 2*XL
J1 IN 0 J(2)
J2 N005260 0 J(2)
J3 N005261 0 J(2)
J4 N005520 0 J(2)
.ENDS
.END
