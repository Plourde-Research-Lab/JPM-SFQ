* source JTL
.SUBCKT SCHEMATIC1  
.ENDS SCHEMATIC1
