*                                               Revised: Thursday, November 15, 2018
* Z:\CHIP-DESIGN\JPM-SFQ\COMPARATOR\ORCAD\COMPARRevision:
*
*
*
*
*
IJPM N00672 0 IJPM*xi
LJPM N00672 0 LJPM*xl
M1 0 LLM(LJPM, LC, M1*xm)
P1 N00256 0 P1
XDCSFQIN N00256 N00081 DCSFQ
XJTL1 N00081 N00085 JTL
XJTL2 N00085 N00089 JTL
XJTL3 N00089 N00372 JTL
I2 N00372 0 I2
LT1 N00372 N00394 L1*xl
J1 N00394 N00434 J(J1*xj)
I1 N00434 0 I1
LQ1 N00434 N00435 LQ1
J2 N00435 N00601 J(J1*xj)
LC N00601 0 LC*xl
LQ2 N00435 N00436 LQ1
J3  N00436 0 J(J1*xj)
LT2 N00434 N00386 L1*xl
XJTL4 N00386 N00224 JTL
XJTL5 N00224 N00228 JTL
R1 N00228 0 R1
.SUBCKT JTL IN OUT
L1 IN N013780 L1*xl
L2 N013780 N014180 L1*xl
L3 N014180 N013980 L1*xl
I1 N014180 0 i1*xi
L4 N013980 OUT L1*xl
J1 N013780 0 J(J1*xj)
J2 N013980 0 J(J1*xj)
.ENDS
.SUBCKT DCSFQ  IN OUT
LJ1 N006000 N006001 L?
LJ2 N006560 0 L?
LJ3 N005480 0 L?
L1 IN N006180 L1
L2 N00480 N005800 L?
L3 N006001 N00480 L?
I2 N00480 0 I?
L4 N005800 N005600 L?
J1 N006000 N006180 JJ
J2 N006001 N006560 JJ
J3 N005800 N005480 JJ
Lq1 N006180 0 L?
XM1 N005600 OUT JTL0
.ENDS
.SUBCKT JTL0  IN OUT
L1 IN N00249 L1*xl
L2 N00249 N003631 L1*xl
L3 N003631 OUT L3*xl
I1 N00249 0 I1*xi
J1 IN 0 J(J1*xj)
J2 N003631 0 J(J1*xj)
.ENDS
.END
