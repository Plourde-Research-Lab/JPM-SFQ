*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision: 
* 
* 
* 
* 
* 
RE1 N00554 0 1.0
P1 N00431 0 Pin
P2 N00475 0 Pin
XJTL1 N00516 N00554 JTL
XJTL2 N00475 N00503 JTL
XJTL N00431 N00512 JTL
Xdff N00503 N00512 N00516 DFF
.SUBCKT JTL  IN OUT
L1 IN N00487 1.0
L2 N00487 N00407 1.0
I1 N00407 0 I1
L3 N00407 N00507 1.0
L4 N00507 OUT 1.0
J1 N00487 0 J
J2 N00507 0 J
.ENDS
.SUBCKT DFF  CLK IN OUT
LJ1 CLK N008111 LJ1
L1 IN N006930 L1
L2 N006930 OUT L2
Lj2 N007211 0 L?
J1 N008111 N006930 JJ
J2 OUT N007211 JJ
.ENDS
.END
