* spice netlist for coupledballisticJTL
* Inductors
L1     1   2   39.5
* Ports
PL1     1   0
PJ1     2   3  2
.end
