*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
RE1 N00554 0 1.0
P1 N00431 0 P1
XJTLIN N00431 N00512 JTL
PCLK N00475 0 PCLK
XJTLCLK N00475 N00503 JTL
XJTLOUT N00516 N00554 JTL
XDFF N00503 N00512 N00516 DFF
.SUBCKT JTL IN OUT
L1 IN N00487 1.0
L2 N00487 N00407 1.0
I1 N00407 0 I1
L3 N00407 N00507 1.0
L4 N00507 OUT 1.0
J1 N00487 0 J
J2 N00507 0 J
.ENDS
.SUBCKT DFF  CLK IN OUT
LJ1 CLK N008111 LJ1
L1 IN N006930 L1
L2 N006930 OUT L2
Lj2 N007211 0 LJ2
J1 N008111 N006930 JJ
J2 OUT N007211 JJ
.ENDS
.SUBCKT SPL1  1 2 3
L1 N020660 N01976 L1*XL
L2 N01976 N021021 L1*XL
I1 N01976 0 I1*XI
L3 3 N01976 L1*XL
L4 1 N020660 L2*XL
L5 N021021 2 L2*XL
J1 N020660 0 JJ
J2 N021021 0 JJ
J3 3 0 JJ
.ENDS
.END
