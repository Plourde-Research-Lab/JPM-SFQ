*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
P1 N00284 0 P1
XDCSFQ N00284 N00214 DCSFQ
XSPL N00214 N00143 N00168 SPL1
RE1 N00143 0 1
RE2 N00168 0 1
.SUBCKT DCSFQ IN OUT
L1 IN N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
Lj1 N004530 N005070 L?
Lj2 N005071 0 L?
Lj3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 OUT JTL1
.ENDS
.SUBCKT JTL1 IN OUT
L1 IN N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 OUT L3*xl
J1 IN 0 JJ
J2 N002320 0 JJ
.ENDS
.SUBCKT SPL1 IN OUT1 OUT2
L1 N020660 N01976 L1*XL
L2 N01976 N021021 L1*XL
I1 N01976 0 I1*XI
L3 IN N01976 L1*XL
L4 OUT1 N020660 L2*XL
L5 N021021 OUT2 L2*XL
J1 N020660 0 JJ
J2 N021021 0 JJ
J3 IN 0 JJ
.ENDS
