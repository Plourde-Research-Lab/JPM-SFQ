* spice netlist 
* Inductors
LJPM      1   2   1000
* Ports
P1     1   2
.end
