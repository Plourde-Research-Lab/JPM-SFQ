*                                               Revised: Thursday, September 13, 2018
* Z:\CHIP-DESIGN\SFQ\JPM RACE ARBITER\JPM RACE ARevision:
*
*
*
*
*
LJPM N08420 0 LJPM*xl
JJPM N08420 0 JT(JJPM*xj)
CJPM N08420 0 CJPM*xc
MA 0 LLM(LJPM, LA1, M1*xm)
MB 0 LLM(LJPM, LB1, -1*M1*xm)
M1 0 LLM(LJPM, Lbias, MBias)
PTrig N04232 0 PTrig
Pd N05712 0 Pd
PReset N04382 0 PReset
LA1 N07390 N03910 L1
LA2 N08880 N03884 L1
LJA1 N034311 0 LJ1
LJA2 N036550 0 LJ1
I1 N03884 0 IC*xci
IBias N087410 0 IBias
LBias N087410 0 LBias
LB1 N07724 N08893 L1
LB2 N08908 N03884 L1
JA1 N03910 N034311 JT(J1*xj)
JA2 N03884 N036550 JT(J1*xj)
LJB1 N037220 0 LJ1
LJB2 N037970 0 LJ1
JB1 N08893 N037220 JT(J1*xj)
JB2 N03884 N037970 JT(J1*xj)
XJTLCLK  N03884 N05205 JTL
XDFF N05205 N04036 N05510 DFF
XResetDC N04382 N04386 DCSFQ
XMRG1 N04386 N05811 N07207 MRG
XMRG2 N05866 N05712 N03075 MRG
XJTLDATA   N03884 N04036 JTL
XBTLB1 N03134 N07724 BJTL5
XBTLB2 N08893 N08908 BJTL5
XBTLA1 N03096 N07390 BJTL5
XBTLA2 N03910 N08880 BJTL5
XIN1   N07207 N03096 JTL
XTrigDC N04232 N04182 DCSFQ
XIN2   N03075 N03134 JTL
XSPL N04182 N05811 N05866 SPL
XJTLOUT   N05510 N06096 JTL
* XSFQDC N06096 N06538 SFQDC
* C1 N06538 0 C1
.SUBCKT SFQDC  IN OUT
LJ1 N000971 0 LJ1
LJ2 N001991 N00649 LJ2*xl
LJ3 N003131 0 LJ3*xl
LJ4 N002551 N00637 LJ4*xl
LJ5 N003691 0 LJ5*xl
LJ6 N00628 N00933 LJ6*xl
LJ7 N008471 0 LJ7*xl
R1 N00933 0 R1
L1 N00649 N00628 L1*xl
L2 N00628 N00637 L2*xl
I1 OUT 0 I1
L3 IN N00106 L3*xl
L4 N000521 N00279 L4*xl
L5 N00106 N000521 L5*xl
J1 N00106 N000971 J
J2 N00279 N001991 J
J3 N00649 N003131 J
J4 N00279 N002551 J
J5 N00637 N003691 J
J6 N00933 OUT JT(J6*xj)
J7 OUT N008471 J
.ENDS
.SUBCKT JTL  IN OUT
L1 IN N009641 L1*xl
L2 N009641 N009420 L2*xl
I1 N009420 0 i1*xi
L3 N009420 OUT L2*xl
J1 N009641 0 J(J1*xj)
J2 OUT 0 J(J1*xj)
.ENDS
.SUBCKT DFF  CLK IN OUT
LJ1 CLK N002671 LJ1*xl
L1 IN N00357 L1*xl
L2 N00357 OUT L2*xl
J1 N002671 N00357 JJ
J2 OUT 0 JJ
.ENDS
.SUBCKT BJTL5  IN OUT
XBJTL3 N002261 N002581 BJTL
XBJTL4 N002581 N002861 BJTL
XBJTL5 N002861 OUT BJTL
XBJTL1 IN N000171 BJTL
XBJTL2 N000171 N002261 BJTL
.ENDS
.SUBCKT BJTL  IN OUT
L1 IN OUT L1
J1 OUT 0 JT(J1*xj)
.ENDS
.SUBCKT DCSFQ  IN OUT
LJ1 N001180 N001181 L?
LJ2 N002971 0 L?
LJ3 N003161 0 L?
L1 IN N000991 L1
L2 N00480 N001611 L?
L3 N001181 N00480 L?
I2 N00480 0 I?
L4 N001611 N001791 L?
J1 N001180 N000991 JJ
J2 N001181 N002971 JJ
J3 N001611 N003161 JJ
Lq1 N000991 0 L?
XM1 N001791 OUT JTL0
.ENDS
.SUBCKT JTL0  IN OUT
L1 IN N00249 L1*xl
L2 N00249 N000611 L1*xl
L3 N000611 OUT L3*xl
I1 N00249 0 I1*xi
J1 IN 0 J(J1*xj)
J2 N000611 0 J(J1*xj)
.ENDS
.SUBCKT MRG  IN1 IN2 OUT
LP1 0 N003310 LP1*xl
LP2 N001921 N004441 LP2*xl
LP3 N006270 N00663 LP3*xl
LP4 N00600 N00663 LP4*xl
LP5 N004630 N002631 LP5*xl
LP6 N003891 0 LP6*xl
LP7 N003611 0 LP7*xl
I1 N006270 0 I1*xi
LT1 IN1 N001921 LT1*xl
LT2 N002970 OUT LT2*xl
LT3 N00663 N002970 LT3*xl
LT4 IN2 N002631 LT4*xl
J1 N003310 N001921 J(J1*xj)
J2 N004441 N00600 J(J2*xj)
J3 N00600 N004630 J(J3*xj)
J4 N002970 N003891 J(J4*xj)
J5 N002631 N003611 J(J5*xj)
.ENDS
.SUBCKT SPL  IN OUT1 OUT2
L1 N00451 N00647 L1*xl
L2 N00451 N00664 L1*xl
I1 N00451 0 I1*xi
L3 IN N00451 L1*xl
L4 N00647 OUT1 L2*xl
L5 N00664 OUT2 L2*xl
J1 N00647 0 JJ
J2 N00664 0 JJ
J3 IN 0 JJ
.ENDS
.END
