*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
P1 N00284 0 P1
XSFQDC N00284 N00214 SFQDC
RE1 N00214 0 RE1
C1 N00214 0 C1
.SUBCKT SFQDC IN OUT
J1 6 7 J(J1*xj)
J2 3 8 J(J2*xj)
J3 10 13 J(J3*xj)
J4 3 9 J(J4*xj)
J5 11 14 J(J5*xj)
J6 4 OUT JT(J6*xj)
J7 OUT 15 J(J7*xj)
I1 0 5 I1
I2 0 OUT I2
L1 10 12 L1
L2 12 11 L2
L3 IN 6 L3
L4 5 3 L4
L5 6 5 L5
LJ1 7 0 LJ1
LJ2 8 10 LJ2
LJ3 13 0 LJ3
LJ4 9 11 LJ4
LJ5 14 0 LJ5
LJ6 4 12 LJ6
LJ7 15 0 LJ7
R1 4 0 R1
.ENDS
.SUBCKT JTL1 IN OUT
L1 IN N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 OUT L3*xl
J1 IN 0 JJ
J2 N002320 0 JJ
.ENDS
