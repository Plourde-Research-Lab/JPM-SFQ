*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
* IJPM 70 0 IJPM
R 70 0 0.01
LJPM 70 0 LJPM
*
PTrig N01 0 PTrig
XTrigDC N01 1 DCSFQ
XSPL 1 101 201 SPL1
*
PReset 2 0 PReset
XResetDC 2 22 DCSFQ
XMRG1 101 22 1001 MRG
XIN1 1001 102 fjtl
XBTLA1 102 3 PTL5
L1 3 4 L1*xl
J1 4 0 JT(J1*xj)
XBTLA2 4 55 PTL5
XBTLA3 55 5 PTL5
L2 5 6 L1*xl
I1 6 0 IC*xci
J2 6 0 JT(J1*xj)
XJTLCLK 6 7 fjtl
*
Pd 200 0 Pd
XMRG2 201 200 2001 MRG
XIN2 2001 202 fjtl
XBTL3 202 23 PTL5
L3 23 24 L1*xl
J3 24 0 JT(J1*xj)
XBTL4 24 205 PTL5
XBTL42 205 25 PTL5
L4 25 26 L1*xl
I3 26 0 IC*xci
J4 26 0 JT(J1*xj)
XJTLDATA 26 27 fjtl
*
M1 0 llm(LJPM, L1, M1*xm)
M2 0 llm(LJPM, L3, -1*M1*xm)
*
XDFF 27 7 9 dff
XJTLOUT 9 10 fjtl
* XSFQDC 10 11 sfqdc
* Cout 11 0 C1
*
.SUBCKT DCSFQ IN OUT
L1 IN N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
LJ1 N004530 N005070 L?
LJ2 N005071 0 L?
LJ3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 OUT JTL0
.ENDS
.SUBCKT JTL0 IN OUT
L1 IN N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 OUT L3*xl
J1 IN 0 J(J1*xj)
J2 N002320 0 J(J1*xj)
.ENDS
.SUBCKT SPL1 IN OUT1 OUT2
L1 N020660 N01976 L1*XL
L2 N01976 N021021 L1*XL
I1 N01976 0 I1*XI
L3 IN N01976 L1*XL
L4 OUT1 N020660 L2*XL
L5 N021021 OUT2 L2*XL
J1 N020660 0 JJ
J2 N021021 0 JJ
J3 IN 0 JJ
.ENDS
.subckt dff IN CLK OUT
LJ1 CLK N008111 LJ1*xl
L1 IN N006930 L1*xl
L2 N006930 OUT L2*xl
Lj2 N007211 0 LJ2*xl
J1 N008111 N006930 JJ
J2 OUT N007211 JJ
.ends dff
.subckt sfqdc IN OUT
J1 6 7 J
J2 3 8 J
J3 10 13 J
J4 3 9 J
J5 11 14 J
J6 4 OUT JT(J6*xj)
J7 OUT 15 J
I1 0 5 I1
I2 0 OUT I2
L1 10 12 L1
L2 12 11 L2
L3 IN 6 L3
L4 5 3 L4
L5 6 5 L5
LJ1 7 0 LJ1
LJ2 8 10 LJ2
LJ3 13 0 LJ3
LJ4 9 11 LJ4
LJ5 14 0 LJ5
LJ6 4 12 LJ6
LJ7 15 0 LJ7
R1 4 0 R1
.ends sfqdc
.subckt fjtl IN OUT
L1 IN 1 L1
J1 1 0 J(J1*xj)
L2 1 2 L2
I1 0 2 I1
L3 2 OUT L2
J2 OUT 0 J(J1*xj)
.ends fjtl
.subckt PTL5 IN OUT
L0 IN 3 L1
J0 3 0 JT(J1*xj)
L1 3 4 L1
J1 4 0 JT(J1*xj)
L2 4 5 L1
J2 5 0 JT(J1*xj)
L3 5 6 L1
J3 6 0 JT(J1*xj)
L4 6 OUT L1
J4 OUT 0 JT(J1*xj)
.ends PTL5
.SUBCKT MRG IN1 IN2 OUT
J1 6 5 J(J1*xj)
J2 4 7 J(J2*xj)
J3 4 11 J(J3*xj)
J4 10 12 J(J4*xj)
J5 13 14 J(J5*xj)
I1 0 8 I1*xi
LP1 0 5 LP1*xl
LP2 7 6 LP2*xl
LP3 8 9 LP3*xl
LP4 4 9 LP4*xl
LP5 11 13 LP5*xl
LP6 0 12 LP6*xl
LP7 0 14 LP7*xl
LT1 IN1 6 LT1*xl
LT2 10 OUT LT2*xl
LT3 9 10 LT3*xl
LT4 IN2 13 LT4*xl
.ENDS
.END
