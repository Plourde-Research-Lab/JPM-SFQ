* spice netlist for InductEx4
L1     1   2   50
L2     3   4   50
L3     5   6   50
* Ports
PL1     1   0
PL2     3   0
PL3     5   0
J1      7   0   10
J2      8   0   10
J3      9   0   10
* JBias   10   0   22.5
.end
