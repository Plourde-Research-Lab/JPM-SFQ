*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
RE1 N00554 0 1.0
P1 N00431 0 P1
XIN N00431 N00432 STDIN
XJTLIN N00431 N00512 JTL1
PCLK N00475 0 PCLK
XCLK N00475 N00476 STDIN
XJTLCLK N00476 N00503 JTL1
XDFF N00503 N00512 N00516 DFF
XJTLOUT N00516 N00554 JTL
XOUT N00554 stdout
.SUBCKT STDIN IN OUT
L1 IN N00519 2*xl
XM1 N00519 N00499 JTL0
XM2 N00499 OUT JTL0
.ENDS
.SUBCKT JTL0 IN OUT
L1 IN N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 OUT L3*xl
J1 IN 0 J(J1*xj)
J2 N002320 0 J(J1*xj)
.ENDS
.SUBCKT JTL1 IN OUT
L1 IN N00487 L1*xl
L2 N00487 N00407 L2*xl
I1 N00407 0 I1*xi
L3 N00407 OUT L2*xl
J1 N00487 0 J(J1*xj)
J2 OUT 0 J(J1*xj)
.ENDS
.SUBCKT JTL IN OUT
L1 IN N00487 L1*xl
L2 N00487 N00407 L2*xl
I1 N00407 0 I1*xi
L3 N00407 N00507 L2*xl
L4 N00507 OUT L1*xl
J1 N00487 0 J(J1*xj)
J2 N00507 0 J(J1*xj)
.ENDS
.SUBCKT DFF  CLK IN OUT
LJ1 CLK N008111 LJ1*xl
L1 IN N006930 L1*xl
L2 N006930 OUT L2*xl
Lj2 N007211 0 LJ2*xl
J1 N008111 N006930 JJ
J2 OUT N007211 JJ
.ENDS
.SUBCKT stdout  IN
R1 N006161 0 0.5
L2 IN N006421 0.75*XL
L3 N006421 N005260 0.75*XL
I1 N006421 0 2.8*XI
L4 N005260 N005261 1.5*XL
I2 N005700 0 2.8*XI
L5 N005261 N005700 0.75*XL
L6 N005700 N005520 0.75*XL
L7 N005520 N006161 2*XL
J1 IN 0 J(2)
J2 N005260 0 J(2)
J3 N005261 0 J(2)
J4 N005520 0 J(2)
.ENDS
.END
