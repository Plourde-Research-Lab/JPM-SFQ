*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
P1 N00284 0 P1
IJPM N005330 0 IJPM
LJPM N005330 0 LJPM
JB1 N00700 0 JT(JB1)
L3 N00700 N00696 L1*XL
JB2 N00692 0 JT(JB2)
L2 N00688 N00692 L1*XL
XDCSFQ N00284 N00214 DCSFQ
XSPL N00214 N00143 N00168 SPL1
XBJTL5 N00143 N00688 BJTL5
XBJTL6 N00692 N00326 BJTL5
XBJTL7 N00180 N00696 BJTL5
XBJTL8 N00700 N00335 BJTL5
XMJTLCLK N00326 N00188 JTL
XMTFF N00168 N00180 TFF
XMJTLIN N00335 N00339 JTL
XJTLOUT N00372 N00376 JTL
XDFF N00188 N00339 N00372 DFF
RE1 N00376 0 1
.SUBCKT JTL IN OUT
L1 IN N00487 1.0
L2 N00487 N00407 1.0
I1 N00407 0 I1
L3 N00407 N00507 1.0
L4 N00507 OUT 1.0
J1 N00487 0 JJ
J2 N00507 0 JJ
.ENDS
.SUBCKT DFF CLK IN OUT
LJ1 CLK N008111 LJ1
L1 IN N006930 L1
L2 N006930 OUT L2
Lj2 N007211 0 LJ2
J1 N008111 N006930 JJ
J2 OUT N007211 JJ
.ENDS
.SUBCKT SPL1  1 2 3
L1 N020660 N01976 L1*XL
L2 N01976 N021021 L1*XL
I1 N01976 0 I1*XI
L3 3 N01976 L1*XL
L4 1 N020660 L2*XL
L5 N021021 2 L2*XL
J1 N020660 0 JJ
J2 N021021 0 JJ
J3 3 0 JJ
.ENDS
.SUBCKT TFF IN OUT
LJ2 N001321 N00332 LJ2
LJ3 N001641 0 LJ3
LJ5 N001801 0 LJ5
LJ4 N001481 N00316 LJ4
L1 N00332 N00475 L1
L2 N00475 2 L2
I1 N000521 0 I1
L3 1 N000361 L3
L4 N000521 N00336 L4
L5 N000361 N000521 L5
J1 N000361 0 JJ
J2 N00336 N001321 JJ
J3 N00332 N001641 JJ
J4 N00336 N001481 JJ
J5 N00316 N001801 JJ
Lq1 N00475 N00316 Lq1
.ENDS
.SUBCKT DCSFQ OUT IN
L1 IN N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
Lj1 N004530 N005070 L?
Lj2 N005071 0 L?
Lj3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 OUT JTL1
.ENDS
.SUBCKT JTL1 IN OUT
L1 1 N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 2 L3*xl
J1 1 0 JJ
J2 N002320 0 JJ
.ENDS
.SUBCKT BJTL IN OUT
L1 IN OUT L?
J1 OUT 0 JT(J1)
.ENDS
.SUBCKT BJTL5 IN OUT
XBJTL1 IN N1 BJTL
XBJTL2 N1 N2 BJTL
XBJTL3 N2 N3 BJTL
XBJTL4 N3 N4 BJTL
XBJTL5 N4 OUT BJTL
.ENDS
.END
