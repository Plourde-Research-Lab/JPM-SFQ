* spice netlist for InductEx4 user manual example 5
* Inductors
LSpiral     1   2   
* Ports
P1     1   2
.end
