* spice netlist for InductEx4 user manual example 5
* Inductors
L1     1   0   5
* Ports
P1     1   0
.end
