*                                               Revised: Monday, November 26, 2018
* Z:\CHIP-DESIGN\JPM-SFQ\COMPARATORV2\ORCAD\COMPRevision: 
* 
* 
* 
* 
* 
JT N07002 N06870 J1
IJPM N06770 0 IJPM
LIN N06998 N07002 L1
LOUT N06870 N07014 L1
IB1 N06870 0 IB1
IB2 N06998 0 IB2
R1 N07022 0 R1
LJPM N06770 0 LJPM
LC N06826 0 LC
P1 N06978 0 P
JB 0 N06870 J1
JE1 N07268 N06998 J1
JE2 N07268 0 J1
JQ N06826 N06870 J2
XJTL1 N06982 N06986 JTL
XJTL2 N06986 N06990 JTL
XJTL3 N06990 N07268 JTL
XJTL4 N07014 N07018 JTL
XJTL5 N07018 N07022 JTL
XDCSFQIN N06978 N06982 DCSFQ
.SUBCKT JTL  IN OUT
L1 IN N013900 L1*xl
L2 N013900 N014300 L2*xl
L3 N014300 N014100 L2*xl
I1 N014300 0 i1*xi
L4 N014100 OUT L1*xl
J1 N013900 0 J(J1*xj)
J2 N014100 0 J(J1*xj)
.ENDS
.SUBCKT DCSFQ  IN OUT
LJ1 N007280 N007880 L?
LJ2 N008261 0 L?
LJ3 N008060 0 L?
L1 IN N007281 L1
L2 N00480 N007680 L?
L3 N007880 N00480 L?
I2 N00480 0 I?
L4 N007680 N007681 L?
J1 N007280 N007281 JJ
J2 N007880 N008261 JJ
J3 N007680 N008060 JJ
Lq1 N007281 0 L?
XM1 N007681 OUT JTL0
.ENDS
.SUBCKT JTL0  IN OUT
L1 IN N00249 L1*xl
L2 N00249 N003751 L1*xl
L3 N003751 OUT L3*xl
I1 N00249 0 I1*xi
J1 IN 0 J(J1*xj)
J2 N003751 0 J(J1*xj)
.ENDS
.END
