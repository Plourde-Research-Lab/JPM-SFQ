*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
P1 N00168 0 P1
XIN1 N00168 N00214 STDIN
XTL21 N00214 N00217 BJTL5
XBTL1 N00217 N00218 JTL1
XBTL2 N00218 N00219 JTL2
R1 N00219 0 R
P2 N60168 0 P2
XIN2 N60168 N61214 STDIN
XTL23 N61214 N10217 BJTL5
XBTL21 N10217 N10218 JTL1
XBTL22 N10218 N10219 JTL2
R2 N10219 0 R
* XDFF N10219 N00219 N20219 DFF
* XOUT N20219 STDOUT
.SUBCKT STDIN IN OUT
L1 IN N00519 2
XM1 N00519 N00499 JTL0
XM2 N00499 OUT JTL0
.ENDS
.SUBCKT JTL0 IN OUT
L1 IN N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 OUT L3*xl
J1 IN 0 J(J1*xj)
J2 N002320 0 J(J1*xj)
.ENDS
.SUBCKT JTL1 IN OUT
L1 IN N002521 L1*xl
J1 N002521 0 J(J1*xj)
L2 N002521 N003521 L1
L3 N003521 N002320 L1*xl
I1 N003521 0 I1*xi
L4 N002320 OUT L1*xl
J2 N002320 0 J(J1*xj)
.ENDS
* .SUBCKT JTL2 IN OUT
* L1 IN N002521 L1*xl
* J1 N002521 0 J(J1)
* L2 N002521 N003521 L1
* L3 N003521 N002320 L1*xl
* I1 N003521 0 I1*xi
* L4 N002320 OUT L1*xl
* J2 N002320 0 J(J1)
* .ENDS
.SUBCKT JTL2 IN OUT
L1 IN N002521 L1*xl
J1 N002521 0 J(J1*xj)
L2 N002521 N003521 L1*xl
L3 N003521 OUT L1*xl
I1 N003521 0 I1*xi
J2 OUT 0 J(J1*xj)
.ENDS
.SUBCKT BJTL5 IN OUT
L1 IN N1 L1*xl
J1 N1 0 JT(J1*xj)
L2 N1 N2 L1*xl
J2 N2 0 JT(J1*xj)
L3 N2 N3 L1*xl
J3 N3 0 JT(J1*xj)
L4 N3 OUT L1*xl
J4 OUT 0 JT(J1*xj)
* L5 N4 OUT L1*xl
* J5 OUT 0 JT(J1*xj)
.ENDS
.END
