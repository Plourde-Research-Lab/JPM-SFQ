WRspice jj I-V curve demo
*
* One can plot a pretty decent iv curve using transient analysis.
* This will show the differences between the various model options.
*
b1 1 0 jj1 control=v2
v1 2 0 pwl(0 0 2n 70m 4n 0 5n 0)
r1 2 1 100
*
* for rtype=4, vary v2 between 0 and 1 for no gap to full gap
v2 3 0 .5
*
r2 3 0 1
*
* It is interesting to set rtype and delv to different values, and note
* the changes.
*
*Nb 1000 A/cm2   area = 30 square microns
.model jj1 jj(rtype=4,cct=1,icon=10m,vg=2.8m,delv=.1m,
+ icrit=0.3m,r0=100,rn=5.4902,cap=1.14195p)
.tran 5p 5n
* type "run", then "plot -b v(1) (-v1#branch)"
.end
