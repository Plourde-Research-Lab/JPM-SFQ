*                                               Revised: Thursday, November 15, 2018
* Z:\CHIP-DESIGN\JPM-SFQ\COMPARATOR\ORCAD\COMPARRevision: 
* 
* 
* 
* 
* 
IJPM N00672 0 IJPM
IB1 N00434 0 IB1
IB2 N00372 0 IB2
R1 N00228 0 R1
L1 N00372 N00394 L2
L2 N00434 N00386 L2
LJPM N00672 0 LJPM
LC N00601 0 LC
P1 N00256 0 P
J1 N00394 N00434 J1
J2 N00601 N00434 J1
J3 0 N00434 J1
XJTL1 N00081 N00085 JTL
XJTL2 N00085 N00089 JTL
XJTL3 N00089 N00372 JTL
XJTL4 N00386 N00224 JTL
XJTL5 N00224 N00228 JTL
XDCSFQIN N00256 N00081 DCSFQ
.SUBCKT JTL  IN OUT
L1 IN N013780 L1*xl
L2 N013780 N014180 L2*xl
L3 N014180 N013980 L2*xl
I1 N014180 0 i1*xi
L4 N013980 OUT L1*xl
J1 N013780 0 J(J1*xj)
J2 N013980 0 J(J1*xj)
.ENDS
.SUBCKT DCSFQ  IN OUT
LJ1 N006000 N006001 L?
LJ2 N006560 0 L?
LJ3 N005480 0 L?
L1 IN N006180 L1
L2 N00480 N005800 L?
L3 N006001 N00480 L?
I2 N00480 0 I?
L4 N005800 N005600 L?
J1 N006000 N006180 JJ
J2 N006001 N006560 JJ
J3 N005800 N005480 JJ
Lq1 N006180 0 L?
XM1 N005600 OUT JTL0
.ENDS
.SUBCKT JTL0  IN OUT
L1 IN N00249 L1*xl
L2 N00249 N003631 L1*xl
L3 N003631 OUT L3*xl
I1 N00249 0 I1*xi
J1 IN 0 J(J1*xj)
J2 N003631 0 J(J1*xj)
.ENDS
.END
