i1 n0 0 i1
j1 n0 0 jn(j1)
r1 n0 0 5.0
.END
