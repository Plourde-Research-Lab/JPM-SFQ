* TB01                                          Revised: Monday, March 20, 2017
* G:\ALEX\RF\MON33\V1\DESIGN1.DSN               Revision: 
* 
* 
* 
* 
* 
L1 N34709 N34726 L1*XL1*XL
I1 N00194 0 I1*XI1
RL1 0 N34674 RL1*XRL1
P1 N334471 0 P1
XMDRV1 N00194 0 N00129 DRV01
XM1 N001490  N334471 STDIN1
XM2 N34747 N34726 N34674 N00194 N34709 mon33
XM3 N34747 STDOUT
XMT1 N001490 N00159 JTL1
XMT2 N00159 N00129 JTL1
.SUBCKT STDOUT  1
R1 N248211 0 0.5
L2 N247991 N248211 2.0
XMT1 1 N247991 JTL
.ENDS
.SUBCKT JTL  1 2
L1 1 N003961 L1*xl
L2 N003961 2 L1*xl
I1 N003961 0 i1*xi
J1 1 0 J
J2 2 0 J(J1)
.ENDS
.SUBCKT mon33  1 2 3 4 5
0 0 0 
Lin1 2 3 Lin1
Lin2 4 5 Lin2
L2 N034610 N034210 L?
L3 N034210 N033890 L?
L4 N033890 1 L?
I2 N034210 0 I?
Lj1 N037631 N035010 Lj1
Lj2 N034751 0 Lj2
Lj3 N033891 0 Lj3
M1 0 LLM(Lin1,Lt1,LM1)
M2 0 LLM(Lin2,Lt2,LM1)
J1 N033750 0 JJJ
J2 N034610 N034751 JJJ
J3 N033890 N033891 JJ
Lt1 N035010 N034610 Lm1*alm*0.5
Lt2 N033750 N037631 Lm1*alm*0.5
.ENDS
.SUBCKT STDIN1  1 2
L1 2 N00519 2
XM1 N00519 N00499 JTL1
XM2 N00499 1 JTL1
.ENDS
.SUBCKT JTL1  1 2
L1 1 N002781 L1*xl
L2 N002781 N002921 L1*xl
L3 N002921 2 L3*xl
I1 N002781 0 i1*xi
J1 1 0 J
J2 N002921 0 J(J1)
.ENDS
.SUBCKT JTL1  1 2
L1 1 N002781 L1*xl
L2 N002781 N002921 L1*xl
L3 N002921 2 L3*xl
I1 N002781 0 i1*xi
J1 1 0 J
J2 N002921 0 J(J1)
.ENDS
.SUBCKT DRV01  1 2 3
0 0 0 
L1 1 N35776 L1*XL1*XL
L2 1 N35786 L1*XL2*XL
R6 N025520 0 R1
L3 3 N02122 L3*XL
R7 N025280 0 R1
I1 N02122 0 I1*XI
L4 N02122 N02572 L4*XL
L5 N02576 N02122 L4*XL
L6 N025280 N02572 L6*XL6*XL
L7 N025520 N02576 L6*XL7*XL
MI1 0 llm(L1,L6,LM1*XLM1)
MI2 0 llm(L2, L7, LM1*XLM2)
Lj2 N000661 2 Lj2
J1 N35776 2 JJJ
J2 1 N000661 JJJ
J3 N35786 2 JJJ(J1,XJ3,VJ1)
J4 3 0 JJ
J5 N02572 0 JJJ
J6 N02576 0 JJJ(J5,XJ6,Vj5)
.ENDS
.END
