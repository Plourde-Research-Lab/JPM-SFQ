*                                               Revised: Tuesday, September 04, 2018
* Z:\CHIP-DESIGN\SFQ\JPM MODEL\JPM.DSN          Revision:
*
*
*
*
*
CCR N00977 N00731 CCR*xc
Ibias N02671 0 Ibias
CCIN N01187 N02580 CCIN*xc
LJPM N00731 0 LJPM
RJPM N00731 0 RJPM
RLC N01187 0 RL
CS N00731 0 CS
Lbias N02671 0 Lbias
RLR N00977 0 RL
JJPM N00731 0 JT(JJPM*xj)
CCC N01052 N00731 CCC*xc
XCavity N02580 N01052 CaptureCavity
MBias 0 LLM(LJPM, Lbias, Mbias)
.SUBCKT CaptureCavity  IN OUT
L1 IN N01680 Ll
L2 N01680 N01799 Ll
L3 N01799 N02464 Ll
L4 N02464 N02431 Ll
L5 N02431 N02038 Ll
L6 N02038 N02042 Ll
L7 N02042 N02046 Ll
C1 IN 0 Cl
L8 N02046 N02236 Ll
C2 N01680 0 Cl
L9 N02236 N02240 Ll
C3 N01799 0 Cl
C4 N02464 0 Cl
C5 N02431 0 Cl
C6 N02038 0 Cl
C7 N02042 0 Cl
C8 N02046 0 Cl
C9 N02236 0 Cl
C10 N02240 0 Cl
L10 N02240 OUT Ll
.ENDS
.END
