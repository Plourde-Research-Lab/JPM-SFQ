*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
P1 N0 0 P1
XDCSFQ N1 N0 DCSFQ
XSPL N2 N3 N1 SPL1
XT1 N3 N11 TFF
XJTLIN N11 N00512 JTL
XJTLCLK N2 N00503 JTL
XDFF N00503 N00512 N00516 DFF
XJTLOUT N00516 N00554 JTL
RE1 N00554 0 1.0
.SUBCKT JTL  IN OUT
L1 IN N00487 1.0
L2 N00487 N00407 1.0
I1 N00407 0 I1
L3 N00407 N00507 1.0
L4 N00507 OUT 1.0
J1 N00487 0 J
J2 N00507 0 J
.ENDS
.SUBCKT DFF  CLK IN OUT
LJ1 CLK N008111 LJ1
L1 IN N006930 L1
L2 N006930 OUT L2
Lj2 N007211 0 LJ2
J1 N008111 N006930 JJ
J2 OUT N007211 JJ
.ENDS
.SUBCKT SPL1  1 2 3
L1 N020660 N01976 L1*XL
L2 N01976 N021021 L1*XL
I1 N01976 0 I1*XI
L3 3 N01976 L1*XL
L4 1 N020660 L2*XL
L5 N021021 2 L2*XL
J1 N020660 0 JJ
J2 N021021 0 JJ
J3 3 0 JJ
.ENDS
.SUBCKT TFF 1 2
LJ2 N001321 N00332 LJ2
LJ3 N001641 0 LJ3
LJ5 N001801 0 LJ5
LJ4 N001481 N00316 LJ4
L1 N00332 N00475 L1
L2 N00475 2 L2
I1 N000521 0 I1
L3 1 N000361 L3
L4 N000521 N00336 L4
L5 N000361 N000521 L5
J1 N000361 0 JJ
J2 N00336 N001321 JJ
J3 N00332 N001641 JJ
J4 N00336 N001481 JJ
J5 N00316 N001801 JJ
Lq1 N00475 N00316 Lq1
.ENDS
.SUBCKT dcsfq  1 2
L1 2 N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
Lj1 N004530 N005070 L?
Lj2 N005071 0 L?
Lj3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 1 JTL1
.ENDS
.SUBCKT JTL1  1 2
L1 1 N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 2 L3*xl
J1 1 0 J
J2 N002320 0 J(J1)
.ENDS
.END
