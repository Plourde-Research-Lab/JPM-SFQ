*                                               Revised: Thursday, March 29, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN4.DSN            Revision:
*
*
*
*
*
P1 N00284 0 P1
XDCSFQ N00284 N00214 DCSFQ
XTL1 N00214 N00215 BJTL5
XTL2 N00215 N00216 BJTL5
XTL3 N00216 N00217 BJTL5
XJTL1 N00217 N00218 AJTL
* XOUT N00217 stdout
R1 N00218 0 R1
.SUBCKT DCSFQ IN OUT
L1 IN N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
Lj1 N004530 N005070 L?
Lj2 N005071 0 L?
Lj3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 OUT JTL1
.ENDS
.SUBCKT JTL1 IN OUT
L1 IN N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 I1*xi
L3 N002320 OUT L3*xl
J1 IN 0 JJ
J2 N002320 0 JJ
.ENDS
.SUBCKT BJTL5 IN OUT
L1 IN N1 L1
J1 N1 0 JT(J1)
L2 N1 N2 L1
J2 N2 0 JT(J1)
L3 N2 N3 L1
J3 N3 0 JT(J1)
L4 N3 N4 L1
J4 N4 0 JT(J1)
L5 N4 OUT L1
J5 OUT 0 JT(J1)
.ENDS
.SUBCKT AJTL IN OUT
L1 IN N1 L1
J1 N1 0 J(J1)
L2 N1 N2 L2
J2 OUT 0 J(J2)
I1 N2 0 I1
L3 N2 OUT L3
.ENDS
.SUBCKT stdout  IN
R0 IN 0 R0
R1 N006161 0 R1
L2 IN N006421 L2*XL
L3 N006421 N005260 L3*XL
I1 N006421 0 I1*XI
L4 N005260 N005261 L4*XL
I2 N005700 0 I1*XI
L5 N005261 N005700 L5*XL
L6 N005700 N005520 L6*XL
L7 N005520 N006161 L7*XL
J1 IN 0 J(J1)
J2 N005260 0 J(J1)
J3 N005261 0 J(J1)
J4 N005520 0 J(J1)
.ENDS
