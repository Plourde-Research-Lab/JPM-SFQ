* SFQ Qbit control                              Revised: Wednesday, February 21, 2018
* root                                          Revision: 2
* A.Kirichenko, HYPRES, INC.
*
*
*
*
I1 N056311 0 I1
XM1 N09052 N056311 dcsfq
XM3 N09246 N09134 N09052 SPL1
.SUBCKT SPL1  1 2 3
L1 N020660 N01976 L1*XL
L2 N01976 N021021 L1*XL
I1 N01976 0 I1*XI
L3 3 N01976 L1*XL
L4 1 N020660 L2*XL
L5 N021021 2 L2*XL
J1 N020660 0 JJ
J2 N021021 0 JJ
J3 3 0 JJ
.ENDS
.SUBCKT dcsfq  1 2
L1 2 N004531 0.1
L2 N004930 N004670 L?
L3 N005070 N004930 L?
I2 N004930 0 I?
L4 N004670 N00693 L?
Lj1 N004530 N005070 L?
Lj2 N005071 0 L?
Lj3 N004671 0 L?
J1 N004530 N004531 JJ
J2 N005070 N005071 JJ
J3 N004670 N004671 JJ
Lq1 N004531 0 L?
XM1 N00693 1 JTL1
.ENDS
.SUBCKT JTL1  1 2
L1 1 N002521 L1*xl
L2 N002521 N002320 L1*xl
I1 N002521 0 i1*xi
L3 N002320 2 L3*xl
J1 1 0 J
J2 N002320 0 J(J1)
.ENDS
.END
