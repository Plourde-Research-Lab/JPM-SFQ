*                                               Revised: Thursday, February 15, 2018
* Z:\CHIP-DESIGN\SFQ\JTL\DESIGN1.DSN            Revision: 
* 
* 
* 
* 
* 
0 0 0 
I2 N36086 0 I
P1 N00130 0 P
XMOUT N00466 STDOUT
XMJTL N00450 N00454 N36086 0 MJTL
XNJTL1 N36125 N00442 NJTL
XNJTL2 N00442 N00446 NJTL
XNJTL3 N00446 N00450 NJTL
XNJTL4 N00454 N00458 NJTL
XMIN N36125 N00130 STDIN
XNJTL5 N00458 N00462 NJTL
XNJTL6 N00462 N00466 NJTL
.SUBCKT STDOUT  1
R1 N250491 0 0.5
L1 1 N25073 L1*XL
L2 N25123 N250491 2.0
XMT1 N25073 N25123 JTL
.ENDS
.SUBCKT JTL  1 2
L2 1 N048790 L1*xl
L3 N048790 N049151 L1*xl
L4 N049151 2 L3*xl
I2 N048790 0 i1*xi
J2 1 0 J
J3 N049151 0 J(J1)
.ENDS
.SUBCKT STDIN  1 2
L1 2 N00612 2
XM1 N00612 N00616 JTL
XM2 N00616 1 JTL
.ENDS
.SUBCKT NJTL  1 2
L1 1 2 L1*XL
I1 2 0 I1*XI1*XI
J1 2 0 JJJ
.ENDS
.SUBCKT MJTL  1 2 3 4
0 0 0 
Lin1 3 4 Lin1*XL
L1 1 2 L1*XL
I1 2 0 I1*XI1*XI
M1 0 LLM(Lin1,L1,LM1)
J1 2 0 JJJ
.ENDS
.END
